`ifndef SRAM_DP_HDE_PARAMS
`define SRAM_DP_HDE_PARAMS

`define WORDS      512
`define BITS       32
`define ADDR_WIDTH $clog2(`WORDS)

`endif  // SRAM_DP_HDE_PARAMS