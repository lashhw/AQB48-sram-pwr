`ifndef RF_2P_HSE_PARAMS
`define RF_2P_HSE_PARAMS

`define WORDS      16
`define BITS       64
`define ADDR_WIDTH $clog2(`WORDS)

`endif  // RF_2P_HSE_PARAMS